module winnerA
(
  input logic [2:0] inA,
  input logic [2:0] inB,
  output logic winA
);

  /*
	Code Here
  */
  
endmodule