
module testbench;

logic ;





endmodule
