module testing (A, B);
    
    input A;
    output B;

    assign B = A;

endmodule
