module validIO
(
  input logic [2:0] inA,
  input logic [2:0] inB,
  output logic valid
);

  /*
	Code Here
  */
  
endmodule