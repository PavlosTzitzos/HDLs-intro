module X_ROM (
	input logic [6:0] address,
	output logic [99:0] data
  );
	always_comb begin
		case (address)
			7'b0000000: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0000001: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0000010: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0000011: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0000100: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0000101: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0000110: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0000111: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0001000: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0001001: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0001010: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0001011: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b0001100: data = 100'b1111111111111111111111111000000000000000000000000000000000000000000000000001111111111111111111111111;
      7'b0001101: data = 100'b0111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111110;
      7'b0001110: data = 100'b0011111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111100;
      7'b0001111: data = 100'b0001111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111000;
      7'b0010000: data = 100'b0000111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111110000;
      7'b0010001: data = 100'b0000011111111111111111111111110000000000000000000000000000000000000000111111111111111111111111100000;
      7'b0010010: data = 100'b0000001111111111111111111111111000000000000000000000000000000000000001111111111111111111111111000000;
      7'b0010011: data = 100'b0000000111111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000;
      7'b0010100: data = 100'b0000000011111111111111111111111110000000000000000000000000000000000111111111111111111111111100000000;
      7'b0010101: data = 100'b0000000001111111111111111111111111000000000000000000000000000000001111111111111111111111111000000000;
      7'b0010110: data = 100'b0000000000111111111111111111111111100000000000000000000000000000011111111111111111111111110000000000;
      7'b0010111: data = 100'b0000000000011111111111111111111111110000000000000000000000000000111111111111111111111111100000000000;
      7'b0011000: data = 100'b0000000000001111111111111111111111111000000000000000000000000001111111111111111111111111000000000000;
      7'b0011001: data = 100'b0000000000000111111111111111111111111100000000000000000000000011111111111111111111111110000000000000;
      7'b0011010: data = 100'b0000000000000011111111111111111111111110000000000000000000000111111111111111111111111100000000000000;
      7'b0011011: data = 100'b0000000000000001111111111111111111111111000000000000000000001111111111111111111111111000000000000000;
      7'b0011100: data = 100'b0000000000000000111111111111111111111111100000000000000000011111111111111111111111110000000000000000;
      7'b0011101: data = 100'b0000000000000000011111111111111111111111110000000000000000111111111111111111111111100000000000000000;
      7'b0011110: data = 100'b0000000000000000001111111111111111111111111000000000000001111111111111111111111111000000000000000000;
      7'b0011111: data = 100'b0000000000000000000111111111111111111111111100000000000011111111111111111111111110000000000000000000;
      7'b0100000: data = 100'b0000000000000000000011111111111111111111111110000000000111111111111111111111111100000000000000000000;
      7'b0100001: data = 100'b0000000000000000000001111111111111111111111111000000001111111111111111111111111000000000000000000000;
      7'b0100010: data = 100'b0000000000000000000000111111111111111111111111100000011111111111111111111111110000000000000000000000;
      7'b0100011: data = 100'b0000000000000000000000011111111111111111111111110000111111111111111111111111100000000000000000000000;
      7'b0100100: data = 100'b0000000000000000000000001111111111111111111111111001111111111111111111111111000000000000000000000000;
      7'b0100101: data = 100'b0000000000000000000000000111111111111111111111111111111111111111111111111110000000000000000000000000;
      7'b0100110: data = 100'b0000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000;
      7'b0100111: data = 100'b0000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000;
      7'b0101000: data = 100'b0000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000;
      7'b0101001: data = 100'b0000000000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000000;
      7'b0101010: data = 100'b0000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000;
      7'b0101011: data = 100'b0000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000;
      7'b0101100: data = 100'b0000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000;
      7'b0101101: data = 100'b0000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000;
      7'b0101110: data = 100'b0000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000;
      7'b0101111: data = 100'b0000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000;
      7'b0110000: data = 100'b0000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000;
      7'b0110001: data = 100'b0000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000;
      7'b0110010: data = 100'b0000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000;
      7'b0110011: data = 100'b0000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000;
      7'b0110100: data = 100'b0000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000;
      7'b0110101: data = 100'b0000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000;
      7'b0110110: data = 100'b0000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000;
      7'b0110111: data = 100'b0000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000;
      7'b0111000: data = 100'b0000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000;
      7'b0111001: data = 100'b0000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000;
      7'b0111010: data = 100'b0000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000;
      7'b0111011: data = 100'b0000000000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000000;
      7'b0111100: data = 100'b0000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000;
      7'b0111101: data = 100'b0000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000;
      7'b0111110: data = 100'b0000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000;
      7'b0111111: data = 100'b0000000000000000000000000111111111111111111111111111111111111111111111111110000000000000000000000000;
      7'b1000000: data = 100'b0000000000000000000000001111111111111111111111111001111111111111111111111111000000000000000000000000;
      7'b1000001: data = 100'b0000000000000000000000011111111111111111111111110000111111111111111111111111100000000000000000000000;
      7'b1000010: data = 100'b0000000000000000000000111111111111111111111111100000011111111111111111111111110000000000000000000000;
      7'b1000011: data = 100'b0000000000000000000001111111111111111111111111000000001111111111111111111111111000000000000000000000;
      7'b1000100: data = 100'b0000000000000000000011111111111111111111111110000000000111111111111111111111111100000000000000000000;
      7'b1000101: data = 100'b0000000000000000000111111111111111111111111100000000000011111111111111111111111110000000000000000000;
      7'b1000110: data = 100'b0000000000000000001111111111111111111111111000000000000001111111111111111111111111000000000000000000;
      7'b1000111: data = 100'b0000000000000000011111111111111111111111110000000000000000111111111111111111111111100000000000000000;
      7'b1001000: data = 100'b0000000000000000111111111111111111111111100000000000000000011111111111111111111111110000000000000000;
      7'b1001001: data = 100'b0000000000000001111111111111111111111111000000000000000000001111111111111111111111111000000000000000;
      7'b1001010: data = 100'b0000000000000011111111111111111111111110000000000000000000000111111111111111111111111100000000000000;
      7'b1001011: data = 100'b0000000000000111111111111111111111111100000000000000000000000011111111111111111111111110000000000000;
      7'b1001100: data = 100'b0000000000001111111111111111111111111000000000000000000000000001111111111111111111111111000000000000;
      7'b1001101: data = 100'b0000000000011111111111111111111111110000000000000000000000000000111111111111111111111111100000000000;
      7'b1001110: data = 100'b0000000000111111111111111111111111100000000000000000000000000000011111111111111111111111110000000000;
      7'b1001111: data = 100'b0000000001111111111111111111111111000000000000000000000000000000001111111111111111111111111000000000;
      7'b1010000: data = 100'b0000000011111111111111111111111110000000000000000000000000000000000111111111111111111111111100000000;
      7'b1010001: data = 100'b0000000111111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000;
      7'b1010010: data = 100'b0000001111111111111111111111111000000000000000000000000000000000000001111111111111111111111111000000;
      7'b1010011: data = 100'b0000011111111111111111111111110000000000000000000000000000000000000000111111111111111111111111100000;
      7'b1010100: data = 100'b0000111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111110000;
      7'b1010101: data = 100'b0001111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111000;
      7'b1010110: data = 100'b0011111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111100;
      7'b1010111: data = 100'b0111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111110;
      7'b1011000: data = 100'b1111111111111111111111111000000000000000000000000000000000000000000000000001111111111111111111111111;
      7'b1011001: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1011010: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1011011: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1011100: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1011101: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1011110: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1011111: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1100000: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1100001: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1100010: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      7'b1100011: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      default: data = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		endcase
	end

endmodule









































