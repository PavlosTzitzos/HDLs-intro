module winnerB
(
  input logic [2:0] inA,
  input logic [2:0] inB,
  output logic winB
);

  /*
	Code Here
  */
  
endmodule