module checkTie
(
  input logic [2:0] inA,
  input logic [2:0] inB,
  output logic tie
);

  /*
	Code Here
  */
  
endmodule